library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all;

entity memory_inst is
  port (
    
  );
end entity memory_inst;